LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY InvSBox IS
    PORT (
        input_byte : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        output_byte : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
END ENTITY;

ARCHITECTURE rtl OF InvSBox IS
    TYPE InvSBoxArray IS ARRAY (0 TO 255) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
    CONSTANT InvSBoxLUT : InvSBoxArray := (
        000 => x"52",
        001 => x"09",
        002 => x"6a",
        003 => x"d5",
        004 => x"30",
        005 => x"36",
        006 => x"a5",
        007 => x"38",
        008 => x"bf",
        009 => x"40",
        010 => x"a3",
        011 => x"9e",
        012 => x"81",
        013 => x"f3",
        014 => x"d7",
        015 => x"fb",
        016 => x"7c",
        017 => x"e3",
        018 => x"39",
        019 => x"82",
        020 => x"9b",
        021 => x"2f",
        022 => x"ff",
        023 => x"87",
        024 => x"34",
        025 => x"8e",
        026 => x"43",
        027 => x"44",
        028 => x"c4",
        029 => x"de",
        030 => x"e9",
        031 => x"cb",
        032 => x"54",
        033 => x"7b",
        034 => x"94",
        035 => x"32",
        036 => x"a6",
        037 => x"c2",
        038 => x"23",
        039 => x"3d",
        040 => x"ee",
        041 => x"4c",
        042 => x"95",
        043 => x"0b",
        044 => x"42",
        045 => x"fa",
        046 => x"c3",
        047 => x"4e",
        048 => x"08",
        049 => x"2e",
        050 => x"a1",
        051 => x"66",
        052 => x"28",
        053 => x"d9",
        054 => x"24",
        055 => x"b2",
        056 => x"76",
        057 => x"5b",
        058 => x"a2",
        059 => x"49",
        060 => x"6d",
        061 => x"8b",
        062 => x"d1",
        063 => x"25",
        064 => x"72",
        065 => x"f8",
        066 => x"f6",
        067 => x"64",
        068 => x"86",
        069 => x"68",
        070 => x"98",
        071 => x"16",
        072 => x"d4",
        073 => x"a4",
        074 => x"5c",
        075 => x"cc",
        076 => x"5d",
        077 => x"65",
        078 => x"b6",
        079 => x"92",
        080 => x"6c",
        081 => x"70",
        082 => x"48",
        083 => x"50",
        084 => x"fd",
        085 => x"ed",
        086 => x"b9",
        087 => x"da",
        088 => x"5e",
        089 => x"15",
        090 => x"46",
        091 => x"57",
        092 => x"a7",
        093 => x"8d",
        094 => x"9d",
        095 => x"84",
        096 => x"90",
        097 => x"d8",
        098 => x"ab",
        099 => x"00",
        100 => x"8c",
        101 => x"bc",
        102 => x"d3",
        103 => x"0a",
        104 => x"f7",
        105 => x"e4",
        106 => x"58",
        107 => x"05",
        108 => x"b8",
        109 => x"b3",
        110 => x"45",
        111 => x"06",
        112 => x"d0",
        113 => x"2c",
        114 => x"1e",
        115 => x"8f",
        116 => x"ca",
        117 => x"3f",
        118 => x"0f",
        119 => x"02",
        120 => x"c1",
        121 => x"af",
        122 => x"bd",
        123 => x"03",
        124 => x"01",
        125 => x"13",
        126 => x"8a",
        127 => x"6b",
        128 => x"3a",
        129 => x"91",
        130 => x"11",
        131 => x"41",
        132 => x"4f",
        133 => x"67",
        134 => x"dc",
        135 => x"ea",
        136 => x"97",
        137 => x"f2",
        138 => x"cf",
        139 => x"ce",
        140 => x"f0",
        141 => x"b4",
        142 => x"e6",
        143 => x"73",
        144 => x"96",
        145 => x"ac",
        146 => x"74",
        147 => x"22",
        148 => x"e7",
        149 => x"ad",
        150 => x"35",
        151 => x"85",
        152 => x"e2",
        153 => x"f9",
        154 => x"37",
        155 => x"e8",
        156 => x"1c",
        157 => x"75",
        158 => x"df",
        159 => x"6e",
        160 => x"47",
        161 => x"f1",
        162 => x"1a",
        163 => x"71",
        164 => x"1d",
        165 => x"29",
        166 => x"c5",
        167 => x"89",
        168 => x"6f",
        169 => x"b7",
        170 => x"62",
        171 => x"0e",
        172 => x"aa",
        173 => x"18",
        174 => x"be",
        175 => x"1b",
        176 => x"fc",
        177 => x"56",
        178 => x"3e",
        179 => x"4b",
        180 => x"c6",
        181 => x"d2",
        182 => x"79",
        183 => x"20",
        184 => x"9a",
        185 => x"db",
        186 => x"c0",
        187 => x"fe",
        188 => x"78",
        189 => x"cd",
        190 => x"5a",
        191 => x"f4",
        192 => x"1f",
        193 => x"dd",
        194 => x"a8",
        195 => x"33",
        196 => x"88",
        197 => x"07",
        198 => x"c7",
        199 => x"31",
        200 => x"b1",
        201 => x"12",
        202 => x"10",
        203 => x"59",
        204 => x"27",
        205 => x"80",
        206 => x"ec",
        207 => x"5f",
        208 => x"60",
        209 => x"51",
        210 => x"7f",
        211 => x"a9",
        212 => x"19",
        213 => x"b5",
        214 => x"4a",
        215 => x"0d",
        216 => x"2d",
        217 => x"e5",
        218 => x"7a",
        219 => x"9f",
        220 => x"93",
        221 => x"c9",
        222 => x"9c",
        223 => x"ef",
        224 => x"a0",
        225 => x"e0",
        226 => x"3b",
        227 => x"4d",
        228 => x"ae",
        229 => x"2a",
        230 => x"f5",
        231 => x"b0",
        232 => x"c8",
        233 => x"eb",
        234 => x"bb",
        235 => x"3c",
        236 => x"83",
        237 => x"53",
        238 => x"99",
        239 => x"61",
        240 => x"17",
        241 => x"2b",
        242 => x"04",
        243 => x"7e",
        244 => x"ba",
        245 => x"77",
        246 => x"d6",
        247 => x"26",
        248 => x"e1",
        249 => x"69",
        250 => x"14",
        251 => x"63",
        252 => x"55",
        253 => x"21",
        254 => x"0c",
        255 => x"7d"
    );
BEGIN
    processInvSBoxLUT : PROCESS (input_byte) IS
    BEGIN
        output_byte <= InvSBoxLUT(to_integer(unsigned(input_byte)));
    END PROCESS;
END ARCHITECTURE;