LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY SBox IS
    PORT (
        input_byte : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        output_byte : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
END ENTITY;

ARCHITECTURE rtl OF SBox IS
    TYPE SBoxArray IS ARRAY (0 TO 255) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
    CONSTANT SBoxLUT : SBoxArray := (
        000 => x"63", 001 => x"7c", 002 => x"77", 003 => x"7b",
        004 => x"f2", 005 => x"6b", 006 => x"6f", 007 => x"c5",
        008 => x"30", 009 => x"01", 010 => x"67", 011 => x"2b",
        012 => x"fe", 013 => x"d7", 014 => x"ab", 015 => x"76",
        016 => x"ca", 017 => x"82", 018 => x"c9", 019 => x"7d",
        020 => x"fa", 021 => x"59", 022 => x"47", 023 => x"f0",
        024 => x"ad", 025 => x"d4", 026 => x"a2", 027 => x"af",
        028 => x"9c", 029 => x"a4", 030 => x"72", 031 => x"c0",
        032 => x"b7", 033 => x"fd", 034 => x"93", 035 => x"26",
        036 => x"36", 037 => x"3f", 038 => x"f7", 039 => x"cc",
        040 => x"34", 041 => x"a5", 042 => x"e5", 043 => x"f1",
        044 => x"71", 045 => x"d8", 046 => x"31", 047 => x"15",
        048 => x"04", 049 => x"c7", 050 => x"23", 051 => x"c3",
        052 => x"18", 053 => x"96", 054 => x"05", 055 => x"9a",
        056 => x"07", 057 => x"12", 058 => x"80", 059 => x"e2",
        060 => x"eb", 061 => x"27", 062 => x"b2", 063 => x"75",
        064 => x"09", 065 => x"83", 066 => x"2c", 067 => x"1a",
        068 => x"1b", 069 => x"6e", 070 => x"5a", 071 => x"a0",
        072 => x"52", 073 => x"3b", 074 => x"d6", 075 => x"b3",
        076 => x"29", 077 => x"e3", 078 => x"2f", 079 => x"84",
        080 => x"53", 081 => x"d1", 082 => x"00", 083 => x"ed",
        084 => x"20", 085 => x"fc", 086 => x"b1", 087 => x"5b",
        088 => x"6a", 089 => x"cb", 090 => x"be", 091 => x"39",
        092 => x"4a", 093 => x"4c", 094 => x"58", 095 => x"cf",
        096 => x"d0", 097 => x"ef", 098 => x"aa", 099 => x"fb",
        100 => x"43", 101 => x"4d", 102 => x"33", 103 => x"85",
        104 => x"45", 105 => x"f9", 106 => x"02", 107 => x"7f",
        108 => x"50", 109 => x"3c", 110 => x"9f", 111 => x"a8",
        112 => x"51", 113 => x"a3", 114 => x"40", 115 => x"8f",
        116 => x"92", 117 => x"9d", 118 => x"38", 119 => x"f5",
        120 => x"bc", 121 => x"b6", 122 => x"da", 123 => x"21",
        124 => x"10", 125 => x"ff", 126 => x"f3", 127 => x"d2",
        128 => x"cd", 129 => x"0c", 130 => x"13", 131 => x"ec",
        132 => x"5f", 133 => x"97", 134 => x"44", 135 => x"17",
        136 => x"c4", 137 => x"a7", 138 => x"7e", 139 => x"3d",
        140 => x"64", 141 => x"5d", 142 => x"19", 143 => x"73",
        144 => x"60", 145 => x"81", 146 => x"4f", 147 => x"dc",
        148 => x"22", 149 => x"2a", 150 => x"90", 151 => x"88",
        152 => x"46", 153 => x"ee", 154 => x"b8", 155 => x"14",
        156 => x"de", 157 => x"5e", 158 => x"0b", 159 => x"db",
        160 => x"e0", 161 => x"32", 162 => x"3a", 163 => x"0a",
        164 => x"49", 165 => x"06", 166 => x"24", 167 => x"5c",
        168 => x"c2", 169 => x"d3", 170 => x"ac", 171 => x"62",
        172 => x"91", 173 => x"95", 174 => x"e4", 175 => x"79",
        176 => x"e7", 177 => x"c8", 178 => x"37", 179 => x"6d",
        180 => x"8d", 181 => x"d5", 182 => x"4e", 183 => x"a9",
        184 => x"6c", 185 => x"56", 186 => x"f4", 187 => x"ea",
        188 => x"65", 189 => x"7a", 190 => x"ae", 191 => x"08",
        192 => x"ba", 193 => x"78", 194 => x"25", 195 => x"2e",
        196 => x"1c", 197 => x"a6", 198 => x"b4", 199 => x"c6",
        200 => x"e8", 201 => x"dd", 202 => x"74", 203 => x"1f",
        204 => x"4b", 205 => x"bd", 206 => x"8b", 207 => x"8a",
        208 => x"70", 209 => x"3e", 210 => x"b5", 211 => x"66",
        212 => x"48", 213 => x"03", 214 => x"f6", 215 => x"0e",
        216 => x"61", 217 => x"35", 218 => x"57", 219 => x"b9",
        220 => x"86", 221 => x"c1", 222 => x"1d", 223 => x"9e",
        224 => x"e1", 225 => x"f8", 226 => x"98", 227 => x"11",
        228 => x"69", 229 => x"d9", 230 => x"8e", 231 => x"94",
        232 => x"9b", 233 => x"1e", 234 => x"87", 235 => x"e9",
        236 => x"ce", 237 => x"55", 238 => x"28", 239 => x"df",
        240 => x"8c", 241 => x"a1", 242 => x"89", 243 => x"0d",
        244 => x"bf", 245 => x"e6", 246 => x"42", 247 => x"68",
        248 => x"41", 249 => x"99", 250 => x"2d", 251 => x"0f",
        252 => x"b0", 253 => x"54", 254 => x"bb", 255 => x"16"
    );
BEGIN
    processSBoxLUT : PROCESS (input_byte) IS
    BEGIN
        output_byte <= SBoxLUT(to_integer(unsigned(input_byte)));
    END PROCESS;
END ARCHITECTURE;